*** SPICE deck for cell tristate_inverter_test{sch} from library Proj2
*** Created on Sun Nov 27, 2016 15:48:52
*** Last revised on Sun Nov 27, 2016 15:52:10
*** Written on Sun Nov 27, 2016 15:53:10 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /home/kenzo/electric/22nm_HP.pm

*** SUBCIRCUIT Proj2__tristate_inverter FROM CELL tristate_inverter{sch}
.SUBCKT Proj2__tristate_inverter EN IN OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 OUT EN net@8 gnd N L=0.022U W=0.176U
Mnmos@2 net@8 IN gnd gnd N L=0.022U W=0.176U
Mnmos@3 net@61 EN gnd gnd N L=0.022U W=0.022U
Mpmos@1 vdd IN net@6 vdd P L=0.022U W=0.176U
Mpmos@2 net@6 net@61 OUT vdd P L=0.022U W=0.176U
Mpmos@3 vdd EN net@61 vdd P L=0.022U W=0.022U
.ENDS Proj2__tristate_inverter

.global gnd vdd

*** TOP LEVEL CELL: tristate_inverter_test{sch}
VVPulse@0 net@3 gnd pulse (0 1V 100ps 200ps 200ps 3ns 6ns) DC 0V AC 0V 0
VVPulse@1 net@7 gnd pulse (0 1V 100ps 200ps 200ps 1.5ns 3ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xtristate@0 net@3 net@7 out Proj2__tristate_inverter
.END
