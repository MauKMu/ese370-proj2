*** SPICE deck for cell bitline_driver{sch} from library Proj2
*** Created on Sat Nov 26, 2016 23:09:06
*** Last revised on Sun Nov 27, 2016 17:39:00
*** Written on Sun Nov 27, 2016 17:39:06 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /home/kenzo/electric/22nm_HP.pm

.global vdd

*** TOP LEVEL CELL: bitline_driver{sch}
Mpmos@0 vdd CLK_ BL_ vdd P L=0.022U W=0.704U
Mpmos@1 vdd CLK_ BL vdd P L=0.022U W=0.704U
.END
