*** SPICE deck for cell d_register_test{sch} from library Proj2
*** Created on Sat Dec 10, 2016 21:56:14
*** Last revised on Sat Dec 10, 2016 22:33:25
*** Written on Sat Dec 10, 2016 22:33:30 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include "C:\Program Files (x86)\Electric\22nm_HP.pm"

*** SUBCIRCUIT Proj2__clk_gen FROM CELL clk_gen{sch}
.SUBCKT Proj2__clk_gen IN OUT OUT_INV
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 A IN gnd gnd N L=0.022U W=0.022U
Mnmos@1 net@3 IN gnd gnd N L=0.022U W=0.022U
Mnmos@2 B net@3 gnd gnd N L=0.022U W=0.022U
Mnmos@3 net@37 A gnd gnd N L=0.022U W=0.022U
Mnmos@4 net@37 OUT_INV gnd gnd N L=0.022U W=0.022U
Mnmos@5 net@50 B gnd gnd N L=0.022U W=0.022U
Mnmos@6 net@50 OUT gnd gnd N L=0.022U W=0.022U
Mnmos@7 net@147 net@37 gnd gnd N L=0.022U W=0.22U
Mnmos@8 OUT net@147 gnd gnd N L=0.022U W=0.022U
Mnmos@9 net@166 net@50 gnd gnd N L=0.022U W=0.22U
Mnmos@10 OUT_INV net@166 gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd IN A vdd P L=0.022U W=0.022U
Mpmos@1 vdd IN net@3 vdd P L=0.022U W=0.022U
Mpmos@2 vdd net@3 B vdd P L=0.022U W=0.022U
Mpmos@3 vdd A net@36 vdd P L=0.022U W=0.022U
Mpmos@4 net@36 OUT_INV net@37 vdd P L=0.022U W=0.022U
Mpmos@5 vdd B net@47 vdd P L=0.022U W=0.022U
Mpmos@6 net@47 OUT net@50 vdd P L=0.022U W=0.022U
Mpmos@7 vdd net@37 net@147 vdd P L=0.022U W=0.22U
Mpmos@8 vdd net@147 OUT vdd P L=0.022U W=0.022U
Mpmos@9 vdd net@50 net@166 vdd P L=0.022U W=0.22U
Mpmos@10 vdd net@166 OUT_INV vdd P L=0.022U W=0.022U
.ENDS Proj2__clk_gen

*** SUBCIRCUIT Proj2__inv FROM CELL inv{sch}
.SUBCKT Proj2__inv x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 y x gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd x y vdd P L=0.022U W=0.022U
.ENDS Proj2__inv

*** SUBCIRCUIT Proj2__nand2 FROM CELL nand2{sch}
.SUBCKT Proj2__nand2 a b y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 y a net@73 gnd N L=0.022U W=0.022U
Mnmos@1 net@73 b gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd a y vdd P L=0.022U W=0.022U
Mpmos@1 vdd b y vdd P L=0.022U W=0.022U
.ENDS Proj2__nand2

*** SUBCIRCUIT Proj2__and2 FROM CELL and2{sch}
.SUBCKT Proj2__and2 a b y
** GLOBAL gnd
** GLOBAL vdd
Xinv@0 net@79 y Proj2__inv
Xnand2@1 a b net@79 Proj2__nand2
.ENDS Proj2__and2

*** SUBCIRCUIT Proj2__nor2 FROM CELL nor2{sch}
.SUBCKT Proj2__nor2 A B Out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Out A gnd gnd N L=0.022U W=0.022U
Mnmos@1 Out B gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A net@0 vdd P L=0.022U W=0.022U
Mpmos@1 net@0 B Out vdd P L=0.022U W=0.022U
.ENDS Proj2__nor2

*** SUBCIRCUIT Proj2__d_latch FROM CELL d_latch{sch}
.SUBCKT Proj2__d_latch In Out φ
** GLOBAL gnd
** GLOBAL vdd
Xand2@0 net@50 φ net@71 Proj2__and2
Xand2@1 φ In net@70 Proj2__and2
Xinv@0 In net@50 Proj2__inv
Xnor2@0 net@71 net@60 Out Proj2__nor2
Xnor2@1 Out net@70 net@60 Proj2__nor2
.ENDS Proj2__d_latch

*** SUBCIRCUIT Proj2__d_register FROM CELL d_register{sch}
.SUBCKT Proj2__d_register D Q φ
** GLOBAL gnd
** GLOBAL vdd
Xclk_gen@1 φ net@31 net@34 Proj2__clk_gen
Xd_latch@2 D net@27 net@34 Proj2__d_latch
Xd_latch@3 net@27 Q net@31 Proj2__d_latch
.ENDS Proj2__d_register

.global gnd vdd

*** TOP LEVEL CELL: d_register_test{sch}
VVPWL@0 D gnd pwl (0ns 0 0.5ns 0 0.5ns 0.8 3.5ns 0.8 3.5ns 0) DC 0V AC 0V 0
VVPulse@0 PHI gnd pulse (0 0.8V 0ns 0 0 1ns 2ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 0.8 AC 0
Xd_regist@0 D Q PHI Proj2__d_register
.END
